interface in_if();
  logic [15:0]a;
  logic [15:0]b;
endinterface
