interface out_if();
  logic [31:0]result;
endinterface
